module unary_not_1_100(A, Z);
    input A;
    output Z;

    assign Z = ~A;
endmodule
