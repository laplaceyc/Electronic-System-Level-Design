module unary_or_2_100(A, Z);
    input [1 : 0] A;
    output Z;

    assign Z = |A;
endmodule
